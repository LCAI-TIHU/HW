module addr_fifo(
    input                   	wclk,
    input                   	rclk,
    input                   	resetn,
    input       [31:0]      	data_in,
    input                   	write_en,
    input                   	read_en,
    output      [31:0]      	data_out,
    output                  	full,
    output                  	empty
);// addr 32
    reg     	[31:0]        	ram[127:0];
    reg     	[7:0]        	write_addr_wclk;
    reg     	[7:0]        	read_addr_rclk;

    wire    	[7:0]        	write_addr_gray_wclk;
    reg     	[7:0]        	write_addr_gray_rclk0;
    reg     	[7:0]        	write_addr_gray_rclk1;

    wire    	[7:0]        	read_addr_gray_rclk;
    reg     	[7:0]        	read_addr_gray_wclk0;
    reg     	[7:0]        	read_addr_gray_wclk1;

    always@(posedge wclk or negedge resetn)//write addr wclk operation
        if(!resetn)
            write_addr_wclk <= 8'b0;
        else if(write_en == 1'b1 && full != 1'b1)
            write_addr_wclk <= write_addr_wclk + 1'b1;
        else
            write_addr_wclk <= write_addr_wclk;
    
    always@(posedge rclk or negedge resetn)//read addr read operation
        if(!resetn)
            read_addr_rclk <= 8'b0;
        else if(read_en == 1'b1 && empty != 1'b1)
            read_addr_rclk <= read_addr_rclk + 1'b1;
        else
            read_addr_rclk <= read_addr_rclk;
    
    always@(posedge wclk or negedge resetn)//sync
        if(!resetn)begin
            read_addr_gray_wclk0 <= 8'b0;
            read_addr_gray_wclk1 <= 8'b0;
        end
        else begin
            read_addr_gray_wclk0 <= read_addr_gray_rclk;
            read_addr_gray_wclk1 <= read_addr_gray_wclk0;
        end
    
    always@(posedge rclk or negedge resetn)//sync
        if(!resetn)begin
            write_addr_gray_rclk0 <= 8'b0;
            write_addr_gray_rclk1 <= 8'b0;
        end
        else begin
            write_addr_gray_rclk0 <= write_addr_gray_wclk;
            write_addr_gray_rclk1 <= write_addr_gray_rclk0;
        end

    always@(posedge wclk or negedge resetn)//data out
		if(!resetn)begin
			ram[0]  <= 31'b0;
			ram[1]  <= 31'b0;
			ram[2]  <= 31'b0;
			ram[3]  <= 31'b0;
			ram[4]  <= 31'b0;
			ram[5]  <= 31'b0;
			ram[6]  <= 31'b0;
			ram[7]  <= 31'b0;
			ram[8]  <= 31'b0;
			ram[9]  <= 31'b0;
			ram[10] <= 31'b0;
			ram[11] <= 31'b0;
			ram[12] <= 31'b0;
			ram[13] <= 31'b0;
			ram[14] <= 31'b0;
			ram[15] <= 31'b0;
			ram[16] <= 31'b0;
			ram[17] <= 31'b0;
			ram[18] <= 31'b0;
			ram[19] <= 31'b0;
			ram[20] <= 31'b0;
			ram[21] <= 31'b0;
			ram[22] <= 31'b0;
			ram[23] <= 31'b0;
			ram[24] <= 31'b0;
			ram[25] <= 31'b0;
			ram[26] <= 31'b0;
			ram[27] <= 31'b0;
			ram[28] <= 31'b0;
			ram[29] <= 31'b0;
			ram[30] <= 31'b0;
			ram[31] <= 31'b0;
			ram[32] <= 31'b0;
			ram[33] <= 31'b0;
			ram[34] <= 31'b0;
			ram[35] <= 31'b0;
			ram[36] <= 31'b0;
			ram[37] <= 31'b0;
			ram[38] <= 31'b0;
			ram[39] <= 31'b0;
			ram[40] <= 31'b0;
			ram[41] <= 31'b0;
			ram[42] <= 31'b0;
			ram[43] <= 31'b0;
			ram[44] <= 31'b0;
			ram[45] <= 31'b0;
			ram[46] <= 31'b0;
			ram[47] <= 31'b0;
			ram[48] <= 31'b0;
			ram[49] <= 31'b0;
			ram[50] <= 31'b0;
			ram[51] <= 31'b0;
			ram[52] <= 31'b0;
			ram[53] <= 31'b0;
			ram[54] <= 31'b0;
			ram[55] <= 31'b0;
			ram[56] <= 31'b0;
			ram[57] <= 31'b0;
			ram[58] <= 31'b0;
			ram[59] <= 31'b0;
			ram[60] <= 31'b0;
			ram[61] <= 31'b0;
			ram[62] <= 31'b0;
			ram[63] <= 31'b0;
			ram[64] <= 31'b0;
			ram[65] <= 31'b0;
			ram[66] <= 31'b0;
			ram[67] <= 31'b0;
			ram[68] <= 31'b0;
			ram[69] <= 31'b0;
			ram[70] <= 31'b0;
			ram[71] <= 31'b0;
			ram[72] <= 31'b0;
			ram[73] <= 31'b0;
			ram[74] <= 31'b0;
			ram[75] <= 31'b0;
			ram[76] <= 31'b0;
			ram[77] <= 31'b0;
			ram[78] <= 31'b0;
			ram[79] <= 31'b0;
			ram[80] <= 31'b0;
			ram[81] <= 31'b0;
			ram[82] <= 31'b0;
			ram[83] <= 31'b0;
			ram[84] <= 31'b0;
			ram[85] <= 31'b0;
			ram[86] <= 31'b0;
			ram[87] <= 31'b0;
			ram[88] <= 31'b0;
			ram[89] <= 31'b0;
			ram[90] <= 31'b0;
			ram[91] <= 31'b0;
			ram[92] <= 31'b0;
			ram[93] <= 31'b0;
			ram[94] <= 31'b0;
			ram[95] <= 31'b0;
			ram[96] <= 31'b0;
			ram[97] <= 31'b0;
			ram[98] <= 31'b0;
			ram[99] <= 31'b0;
			ram[100] <= 31'b0;
			ram[101] <= 31'b0;
			ram[102] <= 31'b0;
			ram[103] <= 31'b0;
			ram[104] <= 31'b0;
			ram[105] <= 31'b0;
			ram[106] <= 31'b0;
			ram[107] <= 31'b0;
			ram[108] <= 31'b0;
			ram[109] <= 31'b0;
			ram[110] <= 31'b0;
			ram[111] <= 31'b0;
			ram[112] <= 31'b0;
			ram[113] <= 31'b0;
			ram[114] <= 31'b0;
			ram[115] <= 31'b0;
			ram[116] <= 31'b0;
			ram[117] <= 31'b0;
			ram[118] <= 31'b0;
			ram[119] <= 31'b0;
			ram[120] <= 31'b0;
			ram[121] <= 31'b0;
			ram[122] <= 31'b0;
			ram[123] <= 31'b0;
			ram[124] <= 31'b0;
			ram[125] <= 31'b0;
			ram[126] <= 31'b0;
			ram[127] <= 31'b0;
		end
        else if(full == 1'b0 && write_en == 1'b1)
            ram[write_addr_wclk[6:0]] <= data_in;


    assign full = (write_addr_gray_wclk[7] != read_addr_gray_wclk1[7])?
                  (write_addr_gray_wclk[6] != read_addr_gray_wclk1[6])?
                  (write_addr_gray_wclk[5:0] == read_addr_gray_wclk1[5:0])?1'b1:1'b0:1'b0:1'b0;
    assign empty = (write_addr_gray_rclk1 == read_addr_gray_rclk)?1'b1:1'b0;
    
	assign data_out = ((read_en == 1'b1) && (empty != 1'b1))?ram[read_addr_rclk[6:0]]:31'b0;
    
	assign write_addr_gray_wclk = (write_addr_wclk>>1)^write_addr_wclk;
    assign read_addr_gray_rclk = (read_addr_rclk>>1)^read_addr_rclk;

endmodule 
